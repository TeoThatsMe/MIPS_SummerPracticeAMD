module Adder(input [31:0] I0,I1,
             output [31:0] out);
  assign out=I0+I1;
endmodule